* /home/ash98/eSim-Workspace/attiny85-test/attiny85-test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat Mar  7 11:58:25 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v2  Net-_U3-Pad1_ GND pulse		
R1  pb0 GND 1k		
U3  Net-_U3-Pad1_ Net-_U3-Pad2_ adc_bridge_1		
U5  Net-_U4-Pad4_ pb0 dac_bridge_1		
U6  pb0 plot_v1		
U1  Net-_U1-Pad1_ GND Net-_U1-Pad3_ Net-_U1-Pad4_ adc_bridge_2		
v1  Net-_U1-Pad1_ GND DC		
U4  Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U3-Pad2_ Net-_U4-Pad4_ ? ? ? ? ? attiny_85_nghdl		

.end
