* /home/shubhangi/eSim-Workspace/exmpl/exmpl.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu Jun 18 18:49:16 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q1  GND Net-_Q1-Pad2_ Net-_Q1-Pad3_ 2N2219		
U3  Net-_U1-Pad4_ Net-_R1-Pad1_ dac_bridge_1		
D1  out3 out4 eSim_LED		
R1  Net-_R1-Pad1_ Net-_Q1-Pad2_ 470		
R3  Net-_Q1-Pad3_ Net-_D3-Pad1_ 150		
R2  out4 Net-_Q1-Pad3_ 150		
U2  out1 GND Net-_U2-Pad3_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ adc_bridge_3		
D3  Net-_D3-Pad1_ out2 eSim_LED		
D4  out2 out1 eSim_LED		
D2  out3 out1 eSim_LED		
v1  out1 GND DC		
v2  Net-_U2-Pad3_ GND pulse		
U5  out3 plot_v1		
U4  out4 plot_v1		
U6  out2 plot_v1		
U7  out1 plot_v1		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ ? ? ? ? ? attiny25		

.end
