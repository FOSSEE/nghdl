
*** input sources ***

v1 100 0 DC PWL ( 0n 0.0 5n 0.0 5.1n 2.0 10n 2.0 10.1n 2.0 15n 2.0 15.1n 0.0 20.0n 0.0 20.1n 2.0 25n 2.0 25.1n 0.0 30n 0.0 30.1n 2.0
		+40.0 2.0 40.1n 0.0 50n 0.0 50.1n 2.0 60n 2.0 60.1n 0.0 70n 0.0 70.1n 2.0 80n 2.0 80.1n 0.0 90n 0.0 100n 0.0)

v2 200 0 DC PWL (0n 2.0 5n 2.0 10n 2.0 15n 2.0 15.1n 0.0 20n 0.0 25n 0.0 30n 0.0 30.1n 2.0 40n 2.0 40.1n 0.0 45n 0.0 45.1n 2.0 
		+ 50n 2.0 50.1n 0.0 60.0n 0.0 70n 0.0 80n 0.0 90n 0.0 95n 0.0 95.1n 2.0 100n 2.0)

Vvdd vdd 0 DC 2.0

*** resistors to ground ***
r1 100 0 1k
r2 200 0 1k


*
*** adc_bridge blocks ***
aconverter1 [100 200 ] [1 2] adc


axor [1] [2]  [12] axors

adac1 [12] [34]  dac
*************model***********

.model axors myxor(rise_delay = 1.0e-10 fall_delay = 1.0e-10 stop_time=90n)

.model adc adc_bridge ( in_low =0.5 in_high =1.0
+                   rise_delay =1.0e-10 fall_delay =1.0e-10)
.model dac dac_bridge(out_low = 0.0 out_high = 2.0 out_undef = 1.0
+                      input_load = 5.0e-14 t_rise = 1.0e-10
+                      t_fall = 1.0e-10)


.end



.CONTROL

option noopalter
tran .1n 100n
.ENDC

