* /home/ash98/eSim-Workspace/piso_test1/piso_test1.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sun Mar 15 16:31:24 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U4  Net-_U1-Pad6_ Serial_Out dac_bridge_1		
R1  Serial_Out GND 1k		
U5  Serial_Out plot_v1		
U3  clock plot_v1		
U1  ? ? ? ? Net-_U1-Pad5_ Net-_U1-Pad6_ piso		
v1  clock GND pulse		
U2  clock Net-_U1-Pad5_ adc_bridge_1		

.end
